module SpaceInvaders (
  input clk,
  input reset, 
  output [7:0] rgb,
  output hSync,
  output vSync,
  );


always @ (clk) begin
 
end     
   

endmodule // SpaceInvaders
